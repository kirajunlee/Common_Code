// ============================================================
// File Name: add_sub_cnt
// VERSION  : V1.0
// DATA     : 2025/02/17
// Author   : lijun
// ============================================================
// 功能：本模块实现计数器加减的操作,支持参数化定义计数器限制的功能;
// ============================================================
module add_sub_cnt #(
    parameter     CNT_WIDTH               = 8                  , //计数器位宽;
    parameter     CNT_LIMIT               = 1'b1                 //计数器限制,即计数器上下溢不做操作;
)
(
    input                                 clk                  ,
    input                                 rst_n                , //复位输入;
    input                                 add                  , //加
    input                                 sub                  , //减
    output logic [CNT_WIDTH-1: 0]         cnt                  , //计数器
    output logic                          cnt_overflow         ,
    output logic                          cnt_underflow
);
//=============================================================
// 本地参数
// ============================================================
//
// ============================================================
// 结构体定义
// ============================================================
//
// ============================================================
// 信号声明
// ============================================================
//
// ============================================================
// 逻辑处理
// ============================================================
always @(posedge clk, negedge rst_n) begin
    if (~rst_n) begin //复位初始化;
        cnt <= 'd0 ;
    end
    else if (add && ~sub) begin //计数器加,但同时没有减操作：
        if ((CNT_LIMIT && ~(&cnt)) || ~CNT_LIMIT) begin //如果计数器限制功能开启,没有计数到最大值计数器才加,或限制关闭只要有加操作计数器就加;
            cnt <= cnt + 1'b1 ;
        end
    end
    else if (~add && sub) begin //计数器减,但同时没有加操作：
        if ((CNT_LIMIT && (|cnt)) || ~CNT_LIMIT) begin //如果计数器限制功能开启,没有计数到0计数器才减,或限制关闭只要有减操作计数器就减 ;
            cnt <= cnt - 1'b1 ;
        end
    end
end

assign cnt_overflow  = (add && ~sub &&  (&cnt))? 1'b1 : 1'b0 ; //加操作但计数器达到最大;
assign cnt_underflow = (~add && sub && ~(|cnt))? 1'b1 : 1'b0 ; //减操作但计数器为0;

endmodule